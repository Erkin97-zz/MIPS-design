module control_unit(opcode, Jump, EX, MEM, WB);
	input [5:0] opcode;

	output reg Jump;
	output reg [3:0] EX; 
	output reg [2:0] MEM; 
	output reg [1:0] WB; 
	
//complete the code
	

endmodule
